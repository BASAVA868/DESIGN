module tb;
 int a;
 initial 
  begin
    $display("test4 folder");
  end

endmodule
